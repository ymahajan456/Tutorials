module hello_world ;

initial begin
  $display ("Hello World by Yogesh");
  #10 $finish;
end

endmodule // End of Module hello_world
